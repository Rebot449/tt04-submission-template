module tt_um_rebot449_lingret_ALU_Top(
    input  wire [7:0] ui_in,    // Dedicated inputs - connected to the input switches
    output wire [7:0] uo_out,   // Dedicated outputs - connected to the 7 segment display
    input  wire [7:0] uio_in,   // IOs: Bidirectional Input path
    output wire [7:0] uio_out,  // IOs: Bidirectional Output path
    output wire [7:0] uio_oe,   // IOs: Bidirectional Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

// use bidirectionals as inputs
    assign uio_oe = 8'b00000000;
// set biderectional output to high impedance
    assign uio_out = 8'bzzzzzzzz;

reg [7:0] r_holder;
always @(ui_in)
begin
	r_holder = ui_in + uio_in;
end
assign uo_out = r_holder;
endmodule
